module	lcd_display_string( 
	clk, 
	rst, 
	index, 
	ones1,
	tens1,
	ones2,
	tens2,
	ones3,
	tens3,
	out);
	
	input				clk;
	input				rst;
	input		[4:0] index;
	input		[3:0]	ones1, tens1, ones2, tens2, ones3, tens3;
	output	[7:0] out;
	
	wire		[3:0]	ones1, tens1, ones2, tens2, ones3, tens3;
	wire		[4:0] index;
	reg		[7:0] out;
	
	always @ ( posedge clk or negedge rst )
		if(!rst)
			out	<=	8'h00;
		else
			case (index)
				00 : out	<=	8'h20;
				01 : out	<=	8'h20;
				02 : out	<=	8'h20;
				03 : out	<=	8'h20;
				04 : out	<=	8'h20;
				05 : out	<=	8'h20;
				06 : out	<=	8'h20;
				07 : out	<=	8'h20;
				08 : out	<=	8'h20;
				09 : out	<=	8'h20;
				10 : out	<=	8'h20;
				11 : out	<=	8'h20;
				12 : out	<=	8'h20;
				13 : out	<=	8'h20;
				14 : out	<=	8'h20;
				15 : out	<=	8'h20;
				
				// line2
				16 : case (tens3)
							0 : out	<=	8'h30;
							1 : out	<= 8'h31;
							2 : out	<= 8'h32;
						default : out <= 8'h20;
					  endcase
				17 : case (ones3)
							0 : out	<=	8'h30;
							1 : out	<= 8'h31;
							2 : out	<= 8'h32;
							3 : out	<= 8'h33;
							4 : out	<= 8'h34;
							5 : out	<= 8'h35;
							6 : out	<= 8'h36;
							7 : out	<= 8'h37;
							8 : out	<= 8'h38;
							9 : out	<= 8'h39;
							default : out <= 8'h20;
					  endcase
				18 : out	<=	8'h3A;
				19 : case (tens2)
							0 : out	<=	8'h30;
							1 : out	<= 8'h31;
							2 : out	<= 8'h32;
							3 : out	<= 8'h33;
							4 : out	<= 8'h34;
							5 : out	<= 8'h35;
						default : out <= 8'h20;
					  endcase
				20 : case (ones2)
							0 : out	<=	8'h30;
							1 : out	<= 8'h31;
							2 : out	<= 8'h32;
							3 : out	<= 8'h33;
							4 : out	<= 8'h34;
							5 : out	<= 8'h35;
							6 : out	<= 8'h36;
							7 : out	<= 8'h37;
							8 : out	<= 8'h38;
							9 : out	<= 8'h39;
							default : out <= 8'h20;
					  endcase
				21 : out	<=	8'h3A;
				22 : case (tens1)
							0 : out	<=	8'h30;
							1 : out	<= 8'h31;
							2 : out	<= 8'h32;
							3 : out	<= 8'h33;
							4 : out	<= 8'h34;
							5 : out	<= 8'h35;
							default : out <= 8'h20;
					  endcase
				23 : case (ones1)
							0 : out	<=	8'h30;
							1 : out	<= 8'h31;
							2 : out	<= 8'h32;
							3 : out	<= 8'h33;
							4 : out	<= 8'h34;
							5 : out	<= 8'h35;
							6 : out	<= 8'h36;
							7 : out	<= 8'h37;
							8 : out	<= 8'h38;
							9 : out	<= 8'h39;
							default : out <= 8'h20;
					  endcase
				24 : out	<=	8'h20;
				25 : out	<=	8'h20;
				26 : out	<=	8'h20;
				27 : out	<=	8'h20;
				28 : out	<=	8'h20;
				29 : out	<=	8'h20;
				30 : out	<=	8'h20;
				31 : out	<=	8'h20;
				default : out <= 8'h20;
			endcase
		
endmodule
				
				
				